----------------------------------------------------------------------------------
-- Company:      TU Wien                                                        --
-- Engineer:     Stefan Adelmann                                                --
--                                                                              --
-- Create Date:  15.03.2018                                                     --
-- Design Name:  Exercise_1                                                     --
-- Module Name:  serial_port_tx_fsm                                             --
-- Project Name: Exercise_1                                                     --
-- Description:  Serial-port transmitter Package                                --
----------------------------------------------------------------------------------

----------------------------------------------------------------------------------
--                                LIBRARIES                                     --
----------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

----------------------------------------------------------------------------------
--                                 PACKAGE                                      --
----------------------------------------------------------------------------------

package serial_port_tx_fsm_pkg is

	--------------------------------------------------------------------
	--                          COMPONENT                             --
	--------------------------------------------------------------------

	-- serial connection of flip-flops to avoid latching of metastable inputs at
	-- the analog/digital interface
	component serial_port_tx_fsm is
		generic (
			CLK_DIVISOR : integer
		);
		port (
			clk : in std_logic;                       --clock
			res_n : in std_logic;                     --low-active reset

			tx : out std_logic;                       --serial output of the parallel input

			data : in std_logic_vector(7 downto 0);   --parallel input byte
			empty : in std_logic;                     --empty signal from the fifo is connected here
			rd : out std_logic                        --connected to the rd input of the fifo
		);
	end component serial_port_tx_fsm;
end package serial_port_tx_fsm_pkg;

--- EOF ---