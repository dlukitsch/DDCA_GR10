library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.core_pack.all;
use work.op_pack.all;

entity ctrl is
	
	port (
            pcsrc : in std_logic;
	    flush_branch : out std_logic
        );

end ctrl;

architecture rtl of ctrl is

begin  -- rtl

    flush_branch <= pcsrc;

end rtl;
